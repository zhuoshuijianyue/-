module top (
    input clk,rst,
    output[7:0] seg0,
    output[7:0] seg1
);
    wire [7:0] f,seg0_not,seg1_not,temp;
    wire f8;
    assign f8=f[7]^f[5]^f[4]^f[3];
    assign temp={f8,f[7:1]};
    Reg #(8, 8'b00010001) u0_reg (clk, rst, temp, f, 1'b1);
   MuxKey #(16, 4, 8) u0_mux (seg0_not, f[3:0], {
    4'd0, 8'b11111100,
    4'd1, 8'b01100000,
    4'd2, 8'b11011010,
    4'd3, 8'b11110010,
    4'd4, 8'b01100110,
    4'd5, 8'b10110110,
    4'd6, 8'b10111110,
    4'd7, 8'b11100000,
    4'd8, 8'b11111110,
    4'd9, 8'b11110110,
    4'd10,8'b11101110,
    4'd11,8'b00111110,
    4'd12,8'b10011100,
    4'd13,8'b01111010,
    4'd14,8'b10011110,
    4'd15,8'b10001110
  });
  MuxKey #(16, 4, 8) u1_mux (seg1_not, f[7:4], {
    4'd0, 8'b11111100,
    4'd1, 8'b01100000,
    4'd2, 8'b11011010,
    4'd3, 8'b11110010,
    4'd4, 8'b01100110,
    4'd5, 8'b10110110,
    4'd6, 8'b10111110,
    4'd7, 8'b11100000,
    4'd8, 8'b11111110,
    4'd9, 8'b11110110,
    4'd10,8'b11101110,
    4'd11,8'b00111110,
    4'd12,8'b10011100,
    4'd13,8'b01111010,
    4'd14,8'b10011110,
    4'd15,8'b10001110
  });
  assign seg0=~seg0_not;
  assign seg1=~seg1_not;
endmodule

